magic
tech sky130A
magscale 1 2
timestamp 1640276982
<< nwell >>
rect 1066 116677 178886 117243
rect 1066 115589 178886 116155
rect 1066 114501 178886 115067
rect 1066 113413 178886 113979
rect 1066 112325 178886 112891
rect 1066 111237 178886 111803
rect 1066 110149 178886 110715
rect 1066 109061 178886 109627
rect 1066 107973 178886 108539
rect 1066 106885 178886 107451
rect 1066 105797 178886 106363
rect 1066 104709 178886 105275
rect 1066 103621 178886 104187
rect 1066 102533 178886 103099
rect 1066 101445 178886 102011
rect 1066 100357 178886 100923
rect 1066 99269 178886 99835
rect 1066 98181 178886 98747
rect 1066 97093 178886 97659
rect 1066 96005 178886 96571
rect 1066 94917 178886 95483
rect 1066 93829 178886 94395
rect 1066 92741 178886 93307
rect 1066 91653 178886 92219
rect 1066 90565 178886 91131
rect 1066 89477 178886 90043
rect 1066 88389 178886 88955
rect 1066 87301 178886 87867
rect 1066 86213 178886 86779
rect 1066 85125 178886 85691
rect 1066 84037 178886 84603
rect 1066 82949 178886 83515
rect 1066 81861 178886 82427
rect 1066 80773 178886 81339
rect 1066 79685 178886 80251
rect 1066 78597 178886 79163
rect 1066 77509 178886 78075
rect 1066 76421 178886 76987
rect 1066 75333 178886 75899
rect 1066 74245 178886 74811
rect 1066 73157 178886 73723
rect 1066 72069 178886 72635
rect 1066 70981 178886 71547
rect 1066 69893 178886 70459
rect 1066 68805 178886 69371
rect 1066 67717 178886 68283
rect 1066 66629 178886 67195
rect 1066 65541 178886 66107
rect 1066 64453 178886 65019
rect 1066 63365 178886 63931
rect 1066 62277 178886 62843
rect 1066 61189 178886 61755
rect 1066 60101 178886 60667
rect 1066 59013 178886 59579
rect 1066 57925 178886 58491
rect 1066 56837 178886 57403
rect 1066 55749 178886 56315
rect 1066 54661 178886 55227
rect 1066 53573 178886 54139
rect 1066 52485 178886 53051
rect 1066 51397 178886 51963
rect 1066 50309 178886 50875
rect 1066 49221 178886 49787
rect 1066 48133 178886 48699
rect 1066 47045 178886 47611
rect 1066 45957 178886 46523
rect 1066 44869 178886 45435
rect 1066 43781 178886 44347
rect 1066 42693 178886 43259
rect 1066 41605 178886 42171
rect 1066 40517 178886 41083
rect 1066 39429 178886 39995
rect 1066 38341 178886 38907
rect 1066 37253 178886 37819
rect 1066 36165 178886 36731
rect 1066 35077 178886 35643
rect 1066 33989 178886 34555
rect 1066 32901 178886 33467
rect 1066 31813 178886 32379
rect 1066 30725 178886 31291
rect 1066 29637 178886 30203
rect 1066 28549 178886 29115
rect 1066 27461 178886 28027
rect 1066 26373 178886 26939
rect 1066 25285 178886 25851
rect 1066 24197 178886 24763
rect 1066 23109 178886 23675
rect 1066 22021 178886 22587
rect 1066 20933 178886 21499
rect 1066 19845 178886 20411
rect 1066 18757 178886 19323
rect 1066 17669 178886 18235
rect 1066 16581 178886 17147
rect 1066 15493 178886 16059
rect 1066 14405 178886 14971
rect 1066 13317 178886 13883
rect 1066 12229 178886 12795
rect 1066 11141 178886 11707
rect 1066 10053 178886 10619
rect 1066 8965 178886 9531
rect 1066 7877 178886 8443
rect 1066 6789 178886 7355
rect 1066 5701 178886 6267
rect 1066 4613 178886 5179
rect 1066 3525 178886 4091
rect 1066 2437 178886 3003
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 2128 178848 117552
<< metal2 >>
rect 2502 0 2558 800
rect 7562 0 7618 800
rect 12714 0 12770 800
rect 17866 0 17922 800
rect 23018 0 23074 800
rect 28170 0 28226 800
rect 33322 0 33378 800
rect 38474 0 38530 800
rect 43626 0 43682 800
rect 48778 0 48834 800
rect 53930 0 53986 800
rect 59082 0 59138 800
rect 64142 0 64198 800
rect 69294 0 69350 800
rect 74446 0 74502 800
rect 79598 0 79654 800
rect 84750 0 84806 800
rect 89902 0 89958 800
rect 95054 0 95110 800
rect 100206 0 100262 800
rect 105358 0 105414 800
rect 110510 0 110566 800
rect 115662 0 115718 800
rect 120814 0 120870 800
rect 125874 0 125930 800
rect 131026 0 131082 800
rect 136178 0 136234 800
rect 141330 0 141386 800
rect 146482 0 146538 800
rect 151634 0 151690 800
rect 156786 0 156842 800
rect 161938 0 161994 800
rect 167090 0 167146 800
rect 172242 0 172298 800
rect 177394 0 177450 800
<< obsm2 >>
rect 2504 856 177448 117552
rect 2614 800 7506 856
rect 7674 800 12658 856
rect 12826 800 17810 856
rect 17978 800 22962 856
rect 23130 800 28114 856
rect 28282 800 33266 856
rect 33434 800 38418 856
rect 38586 800 43570 856
rect 43738 800 48722 856
rect 48890 800 53874 856
rect 54042 800 59026 856
rect 59194 800 64086 856
rect 64254 800 69238 856
rect 69406 800 74390 856
rect 74558 800 79542 856
rect 79710 800 84694 856
rect 84862 800 89846 856
rect 90014 800 94998 856
rect 95166 800 100150 856
rect 100318 800 105302 856
rect 105470 800 110454 856
rect 110622 800 115606 856
rect 115774 800 120758 856
rect 120926 800 125818 856
rect 125986 800 130970 856
rect 131138 800 136122 856
rect 136290 800 141274 856
rect 141442 800 146426 856
rect 146594 800 151578 856
rect 151746 800 156730 856
rect 156898 800 161882 856
rect 162050 800 167034 856
rect 167202 800 172186 856
rect 172354 800 177338 856
<< obsm3 >>
rect 4208 2143 173488 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< labels >>
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 1 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 1 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 1 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 1 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 1 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 1 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 2 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 2 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 2 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 2 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 2 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 2 nsew ground input
rlabel metal2 s 2502 0 2558 800 6 wb_clk_i
port 3 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wb_rst_i
port 4 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_dat_o[0]
port 5 nsew signal output
rlabel metal2 s 69294 0 69350 800 6 wbs_dat_o[10]
port 6 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 wbs_dat_o[11]
port 7 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 wbs_dat_o[12]
port 8 nsew signal output
rlabel metal2 s 84750 0 84806 800 6 wbs_dat_o[13]
port 9 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 wbs_dat_o[14]
port 10 nsew signal output
rlabel metal2 s 95054 0 95110 800 6 wbs_dat_o[15]
port 11 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 wbs_dat_o[16]
port 12 nsew signal output
rlabel metal2 s 105358 0 105414 800 6 wbs_dat_o[17]
port 13 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 wbs_dat_o[18]
port 14 nsew signal output
rlabel metal2 s 115662 0 115718 800 6 wbs_dat_o[19]
port 15 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_o[1]
port 16 nsew signal output
rlabel metal2 s 120814 0 120870 800 6 wbs_dat_o[20]
port 17 nsew signal output
rlabel metal2 s 125874 0 125930 800 6 wbs_dat_o[21]
port 18 nsew signal output
rlabel metal2 s 131026 0 131082 800 6 wbs_dat_o[22]
port 19 nsew signal output
rlabel metal2 s 136178 0 136234 800 6 wbs_dat_o[23]
port 20 nsew signal output
rlabel metal2 s 141330 0 141386 800 6 wbs_dat_o[24]
port 21 nsew signal output
rlabel metal2 s 146482 0 146538 800 6 wbs_dat_o[25]
port 22 nsew signal output
rlabel metal2 s 151634 0 151690 800 6 wbs_dat_o[26]
port 23 nsew signal output
rlabel metal2 s 156786 0 156842 800 6 wbs_dat_o[27]
port 24 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 wbs_dat_o[28]
port 25 nsew signal output
rlabel metal2 s 167090 0 167146 800 6 wbs_dat_o[29]
port 26 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_o[2]
port 27 nsew signal output
rlabel metal2 s 172242 0 172298 800 6 wbs_dat_o[30]
port 28 nsew signal output
rlabel metal2 s 177394 0 177450 800 6 wbs_dat_o[31]
port 29 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_o[3]
port 30 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 wbs_dat_o[4]
port 31 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 wbs_dat_o[5]
port 32 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 wbs_dat_o[6]
port 33 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 wbs_dat_o[7]
port 34 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 wbs_dat_o[8]
port 35 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 wbs_dat_o[9]
port 36 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 wbs_stb_i
port 37 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 5625756
string GDS_START 163558
<< end >>

